6T_SRAM_Read_1
.include "45nm_HP.pm
Vdd d 0 1.1

MM1 Q Qb 0 0 N L=0.05U W=0.1U AS=0.019P AD=0.026P PS=0.575U PD=0.558U
MM2 Q d BL 0 N L=0.05U W=0.15U AS=0.024P AD=0.026P PS=0.625U PD=0.558U
MM3 Q Qb d d P L=0.05U W=0.2U AS=0.033P AD=0.026P PS=0.725U PD=0.558U
MM4 Qb Q 0 0 N L=0.05U W=0.1U AS=0.019P AD=0.026P PS=0.575U PD=0.558U
MM5 BLB d Qb 0 N L=0.05U W=0.15U AS=0.026P AD=0.024P PS=0.558U PD=0.625U
MM6 Qb Q d d P L=0.05U W=0.2U AS=0.033P AD=0.026P PS=0.725U PD=0.558U

Vin1 Q 0 PWL(0ns 0 5ns 0 5.1ns 1.1 10ns 1.1 10.1ns 0 15ns 0 15.1ns 1.1)
Vin2 Qb 0 PWL(0ns 1.1 5ns 1.1 5.1ns 0 10ns 0 10.1ns 1.1 15ns 1.1 15.1ns 0)
.tran 0ps 20ns 0 1ns
.print tran V(Q) V(Qb) V(BL) V(BLB)
.end